* sg13g2_IOPadTriOut24mA
.subckt sg13g2_IOPadTriOut24mA vss vdd iovss iovdd c2p c2p_en pad
Xnclamp iovss iovdd pad ngate sg13g2_Clamp_N12N12D
Xpclamp iovss iovdd pad pgate sg13g2_Clamp_P12N12D
Xdcndiode iovss pad iovdd sg13g2_DCNDiode
Xdcpdiode pad iovdd iovss sg13g2_DCPDiode
Xgatedec vdd vss iovdd c2p c2p_en ngate pgate sg13g2_GateDecode
.ends sg13g2_IOPadTriOut24mA
