* sg13g2_IOPadInOut16mA
.subckt sg13g2_IOPadInOut16mA vss vdd iovss iovdd p2c c2p c2p_en pad
Xnclamp iovss iovdd pad ngate sg13g2_Clamp_N8N8D
Xpclamp iovss iovdd pad pgate sg13g2_Clamp_P8N8D
Xdcndiode iovss pad iovdd sg13g2_DCNDiode
Xdcpdiode pad iovdd iovss sg13g2_DCPDiode
Xgatedec vdd vss iovdd c2p c2p_en ngate pgate sg13g2_GateDecode
Xleveldown vdd vss iovdd iovss pad p2c sg13g2_LevelDown
.ends sg13g2_IOPadInOut16mA
