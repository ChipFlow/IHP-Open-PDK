* sg13g2_Clamp_P20N0D hierarchy

* sg13g2_GuardRing_P16000W3852HFF
.subckt sg13g2_GuardRing_P16000W3852HFF conn

.ends sg13g2_GuardRing_P16000W3852HFF

* sg13g2_GuardRing_N15280W3132HTF
.subckt sg13g2_GuardRing_N15280W3132HTF conn

.ends sg13g2_GuardRing_N15280W3132HTF

* sg13g2_Clamp_P20N0D
.subckt sg13g2_Clamp_P20N0D iovss iovdd pad
Xclamp_g0_r0 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g0_r1 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g1_r0 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g1_r1 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g2_r0 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g2_r1 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g3_r0 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g3_r1 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g4_r0 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g4_r1 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g5_r0 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g5_r1 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g6_r0 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g6_r1 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g7_r0 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g7_r1 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g8_r0 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g8_r1 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g9_r0 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g9_r1 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g10_r0 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g10_r1 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g11_r0 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g11_r1 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g12_r0 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g12_r1 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g13_r0 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g13_r1 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g14_r0 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g14_r1 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g15_r0 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g15_r1 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g16_r0 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g16_r1 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g17_r0 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g17_r1 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g18_r0 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g18_r1 iovdd off pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g19_r0 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g19_r1 pad off iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
XOuterRing iovss sg13g2_GuardRing_P16000W3852HFF
XInnerRing iovdd sg13g2_GuardRing_N15280W3132HTF
RRoff iovdd off 6708.0
.ends sg13g2_Clamp_P20N0D
