* sg13g2_GuardRing_P456W948HFF hierarchy

* sg13g2_GuardRing_P456W948HFF
.subckt sg13g2_GuardRing_P456W948HFF conn

.ends sg13g2_GuardRing_P456W948HFF
