* inv_x1
.subckt inv_x1 vdd vss i nq
Xnmos vss i nq vss sg13_lv_nmos l=0.13um w=3.93um
Xpmos vdd i nq vdd sg13_lv_pmos l=0.13um w=4.41um
.ends inv_x1
