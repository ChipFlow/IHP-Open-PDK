* sg13g2_Filler10000 hierarchy

* sg13g2_Filler10000
.subckt sg13g2_Filler10000 vss vdd iovss iovdd

.ends sg13g2_Filler10000
