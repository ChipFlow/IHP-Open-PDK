* sg13g2_Filler4000 hierarchy

* sg13g2_Filler4000
.subckt sg13g2_Filler4000 vss vdd iovss iovdd

.ends sg13g2_Filler4000
