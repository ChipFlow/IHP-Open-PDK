* sg13g2_Clamp_N43N43D4R hierarchy

* sg13g2_GuardRing_N16000W4884HFF
.subckt sg13g2_GuardRing_N16000W4884HFF conn

.ends sg13g2_GuardRing_N16000W4884HFF

* sg13g2_GuardRing_P15280W4164HFF
.subckt sg13g2_GuardRing_P15280W4164HFF conn

.ends sg13g2_GuardRing_P15280W4164HFF

* sg13g2_Clamp_N43N43D4R
.subckt sg13g2_Clamp_N43N43D4R iovss iovdd pad gate
Xclamp_g0_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g0_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g0_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g0_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g1_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g1_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g1_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g1_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g2_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g2_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g2_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g2_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g3_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g3_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g3_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g3_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g4_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g4_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g4_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g4_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g5_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g5_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g5_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g5_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g6_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g6_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g6_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g6_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g7_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g7_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g7_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g7_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g8_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g8_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g8_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g8_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g9_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g9_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g9_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g9_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g10_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g10_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g10_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g10_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g11_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g11_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g11_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g11_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g12_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g12_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g12_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g12_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g13_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g13_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g13_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g13_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g14_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g14_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g14_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g14_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g15_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g15_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g15_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g15_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g16_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g16_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g16_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g16_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g17_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g17_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g17_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g17_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g18_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g18_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g18_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g18_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g19_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g19_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g19_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g19_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g20_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g20_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g20_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g20_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g21_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g21_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g21_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g21_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g22_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g22_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g22_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g22_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g23_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g23_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g23_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g23_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g24_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g24_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g24_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g24_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g25_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g25_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g25_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g25_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g26_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g26_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g26_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g26_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g27_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g27_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g27_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g27_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g28_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g28_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g28_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g28_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g29_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g29_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g29_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g29_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g30_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g30_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g30_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g30_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g31_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g31_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g31_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g31_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g32_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g32_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g32_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g32_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g33_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g33_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g33_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g33_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g34_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g34_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g34_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g34_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g35_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g35_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g35_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g35_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g36_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g36_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g36_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g36_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g37_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g37_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g37_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g37_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g38_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g38_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g38_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g38_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g39_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g39_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g39_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g39_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g40_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g40_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g40_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g40_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g41_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g41_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g41_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g41_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g42_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g42_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g42_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g42_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
XOuterRing iovdd sg13g2_GuardRing_N16000W4884HFF
XInnerRing iovss sg13g2_GuardRing_P15280W4164HFF
XDGATE iovss gate dantenna l=0.64um w=0.3um
.ends sg13g2_Clamp_N43N43D4R
