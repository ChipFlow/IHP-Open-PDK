* sg13g2_Filler200
.subckt sg13g2_Filler200 vss vdd iovss iovdd

.ends sg13g2_Filler200
