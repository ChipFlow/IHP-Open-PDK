* sg13g2_Filler1000 hierarchy

* sg13g2_Filler1000
.subckt sg13g2_Filler1000 vss vdd iovss iovdd

.ends sg13g2_Filler1000
