* sg13g2_IOPadOut20mA
.subckt sg13g2_IOPadOut20mA vss vdd iovss iovdd c2p pad
Xnclamp iovss iovdd pad ngate sg13g2_Clamp_N10N10D
Xpclamp iovss iovdd pad pgate sg13g2_Clamp_P10N10D
Xdcndiode iovss pad iovdd sg13g2_DCNDiode
Xdcpdiode pad iovdd iovss sg13g2_DCPDiode
Xgatelu vdd vss iovdd c2p ngate pgate sg13g2_GateLevelUpInv
.ends sg13g2_IOPadOut20mA
