* sg13g2_Gallery
.subckt sg13g2_Gallery vdd vss iovdd iopadin_pad iopadout4ma_pad iopadout8ma_pad iopadout12ma_pad iopadout16ma_pad iopadout20ma_pad iopadout24ma_pad iopadout30ma_pad iopadtriout4ma_pad iopadtriout8ma_pad iopadtriout12ma_pad iopadtriout16ma_pad iopadtriout20ma_pad iopadtriout24ma_pad iopadtriout30ma_pad iopadinout4ma_pad iopadinout8ma_pad iopadinout12ma_pad iopadinout16ma_pad iopadinout20ma_pad iopadinout24ma_pad iopadinout30ma_pad iopadin_p2c iopadinout4ma_p2c iopadinout8ma_p2c iopadinout12ma_p2c iopadinout16ma_p2c iopadinout20ma_p2c iopadinout24ma_p2c iopadinout30ma_p2c iopadout4ma_c2p iopadout8ma_c2p iopadout12ma_c2p iopadout16ma_c2p iopadout20ma_c2p iopadout24ma_c2p iopadout30ma_c2p iopadtriout4ma_c2p iopadtriout8ma_c2p iopadtriout12ma_c2p iopadtriout16ma_c2p iopadtriout20ma_c2p iopadtriout24ma_c2p iopadtriout30ma_c2p iopadinout4ma_c2p iopadinout8ma_c2p iopadinout12ma_c2p iopadinout16ma_c2p iopadinout20ma_c2p iopadinout24ma_c2p iopadinout30ma_c2p iopadtriout4ma_c2p_en iopadtriout8ma_c2p_en iopadtriout12ma_c2p_en iopadtriout16ma_c2p_en iopadtriout20ma_c2p_en iopadtriout24ma_c2p_en iopadtriout30ma_c2p_en iopadinout4ma_c2p_en iopadinout8ma_c2p_en iopadinout12ma_c2p_en iopadinout16ma_c2p_en iopadinout20ma_c2p_en iopadinout24ma_c2p_en iopadinout30ma_c2p_en ana_out ana_outres
Xcorner vss vdd vss iovdd sg13g2_Corner
Xfiller200 vss vdd vss iovdd sg13g2_Filler200
Xfiller400 vss vdd vss iovdd sg13g2_Filler400
Xfiller1000 vss vdd vss iovdd sg13g2_Filler1000
Xfiller2000 vss vdd vss iovdd sg13g2_Filler2000
Xfiller4000 vss vdd vss iovdd sg13g2_Filler4000
Xfiller10000 vss vdd vss iovdd sg13g2_Filler10000
Xiopadvss vss vdd vss iovdd sg13g2_IOPadVss
Xiopadvdd vss vdd vss iovdd sg13g2_IOPadVdd
Xiopadin vss vdd vss iovdd iopadin_p2c iopadin_pad sg13g2_IOPadIn
Xiopadout4ma vss vdd vss iovdd iopadout4ma_c2p iopadout4ma_pad sg13g2_IOPadOut4mA
Xiopadout8ma vss vdd vss iovdd iopadout8ma_c2p iopadout8ma_pad sg13g2_IOPadOut8mA
Xiopadout12ma vss vdd vss iovdd iopadout12ma_c2p iopadout12ma_pad sg13g2_IOPadOut12mA
Xiopadout16ma vss vdd vss iovdd iopadout16ma_c2p iopadout16ma_pad sg13g2_IOPadOut16mA
Xiopadout20ma vss vdd vss iovdd iopadout20ma_c2p iopadout20ma_pad sg13g2_IOPadOut20mA
Xiopadout24ma vss vdd vss iovdd iopadout24ma_c2p iopadout24ma_pad sg13g2_IOPadOut24mA
Xiopadout30ma vss vdd vss iovdd iopadout30ma_c2p iopadout30ma_pad sg13g2_IOPadOut30mA
Xiopadtriout4ma vss vdd vss iovdd iopadtriout4ma_c2p iopadtriout4ma_c2p_en iopadtriout4ma_pad sg13g2_IOPadTriOut4mA
Xiopadtriout8ma vss vdd vss iovdd iopadtriout8ma_c2p iopadtriout8ma_c2p_en iopadtriout8ma_pad sg13g2_IOPadTriOut8mA
Xiopadtriout12ma vss vdd vss iovdd iopadtriout12ma_c2p iopadtriout12ma_c2p_en iopadtriout12ma_pad sg13g2_IOPadTriOut12mA
Xiopadtriout16ma vss vdd vss iovdd iopadtriout16ma_c2p iopadtriout16ma_c2p_en iopadtriout16ma_pad sg13g2_IOPadTriOut16mA
Xiopadtriout20ma vss vdd vss iovdd iopadtriout20ma_c2p iopadtriout20ma_c2p_en iopadtriout20ma_pad sg13g2_IOPadTriOut20mA
Xiopadtriout24ma vss vdd vss iovdd iopadtriout24ma_c2p iopadtriout24ma_c2p_en iopadtriout24ma_pad sg13g2_IOPadTriOut24mA
Xiopadtriout30ma vss vdd vss iovdd iopadtriout30ma_c2p iopadtriout30ma_c2p_en iopadtriout30ma_pad sg13g2_IOPadTriOut30mA
Xiopadinout4ma vss vdd vss iovdd iopadinout4ma_p2c iopadinout4ma_c2p iopadinout4ma_c2p_en iopadinout4ma_pad sg13g2_IOPadInOut4mA
Xiopadinout8ma vss vdd vss iovdd iopadinout8ma_p2c iopadinout8ma_c2p iopadinout8ma_c2p_en iopadinout8ma_pad sg13g2_IOPadInOut8mA
Xiopadinout12ma vss vdd vss iovdd iopadinout12ma_p2c iopadinout12ma_c2p iopadinout12ma_c2p_en iopadinout12ma_pad sg13g2_IOPadInOut12mA
Xiopadinout16ma vss vdd vss iovdd iopadinout16ma_p2c iopadinout16ma_c2p iopadinout16ma_c2p_en iopadinout16ma_pad sg13g2_IOPadInOut16mA
Xiopadinout20ma vss vdd vss iovdd iopadinout20ma_p2c iopadinout20ma_c2p iopadinout20ma_c2p_en iopadinout20ma_pad sg13g2_IOPadInOut20mA
Xiopadinout24ma vss vdd vss iovdd iopadinout24ma_p2c iopadinout24ma_c2p iopadinout24ma_c2p_en iopadinout24ma_pad sg13g2_IOPadInOut24mA
Xiopadinout30ma vss vdd vss iovdd iopadinout30ma_p2c iopadinout30ma_c2p iopadinout30ma_c2p_en iopadinout30ma_pad sg13g2_IOPadInOut30mA
Xiopadiovss vss vdd vss iovdd sg13g2_IOPadIOVss
Xiopadiovdd vss vdd vss iovdd sg13g2_IOPadIOVdd
Xiopadanalog vss vdd vss iovdd ana_out ana_outres sg13g2_IOPadAnalog
Xcorner2 vss vdd vss iovdd sg13g2_Corner
.ends sg13g2_Gallery
