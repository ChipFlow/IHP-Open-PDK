* sg13g2_RCClampInverter hierarchy

* sg13g2_GuardRing_P16000W4466HFT
.subckt sg13g2_GuardRing_P16000W4466HFT conn

.ends sg13g2_GuardRing_P16000W4466HFT

* sg13g2_GuardRing_N9472W2216HTT
.subckt sg13g2_GuardRing_N9472W2216HTT conn

.ends sg13g2_GuardRing_N9472W2216HTT

* sg13g2_RCClampInverter
.subckt sg13g2_RCClampInverter supply ground in out
Xcapmos0_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos1_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos2_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos3_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos4_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos5_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos6_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xnmos0_r0 ground in out ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos1_r0 out in ground ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos2_r0 ground in out ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos3_r0 out in ground ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos4_r0 ground in out ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos5_r0 out in ground ground sg13_hv_nmos l=0.5um w=9.0um
Xcapmos0_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos1_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos2_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos3_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos4_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos5_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos6_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xnmos0_r1 ground in out ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos1_r1 out in ground ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos2_r1 ground in out ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos3_r1 out in ground ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos4_r1 ground in out ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos5_r1 out in ground ground sg13_hv_nmos l=0.5um w=9.0um
Xnmosguardring ground sg13g2_GuardRing_P16000W4466HFT
Xpmos0_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos1_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos2_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos3_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos4_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos5_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos6_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos7_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos8_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos9_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos10_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos11_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos12_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos13_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos14_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos15_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos16_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos17_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos18_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos19_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos20_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos21_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos22_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos23_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos24_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos25_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos26_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos27_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos28_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos29_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos30_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos31_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos32_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos33_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos34_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos35_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos36_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos37_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos38_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos39_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos40_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos41_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos42_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos43_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos44_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos45_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos46_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos47_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos48_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos49_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmosguardring supply sg13g2_GuardRing_N9472W2216HTT
.ends sg13g2_RCClampInverter
