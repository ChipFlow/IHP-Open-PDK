* sg13g2_IOPadOut20mA hierarchy

* sg13g2_GuardRing_N16000W1980HFF
.subckt sg13g2_GuardRing_N16000W1980HFF conn

.ends sg13g2_GuardRing_N16000W1980HFF

* sg13g2_GuardRing_P15280W1260HFF
.subckt sg13g2_GuardRing_P15280W1260HFF conn

.ends sg13g2_GuardRing_P15280W1260HFF

* sg13g2_Clamp_N10N10D
.subckt sg13g2_Clamp_N10N10D iovss iovdd pad gate
Xclamp_g0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g4 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g5 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g6 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g7 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g8 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g9 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
XOuterRing iovdd sg13g2_GuardRing_N16000W1980HFF
XInnerRing iovss sg13g2_GuardRing_P15280W1260HFF
XDGATE iovss gate dantenna l=0.64um w=0.3um
.ends sg13g2_Clamp_N10N10D

* sg13g2_GuardRing_P16000W3852HFF
.subckt sg13g2_GuardRing_P16000W3852HFF conn

.ends sg13g2_GuardRing_P16000W3852HFF

* sg13g2_GuardRing_N15280W3132HTF
.subckt sg13g2_GuardRing_N15280W3132HTF conn

.ends sg13g2_GuardRing_N15280W3132HTF

* sg13g2_Clamp_P10N10D
.subckt sg13g2_Clamp_P10N10D iovss iovdd pad gate
Xclamp_g0_r0 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g0_r1 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g1_r0 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g1_r1 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g2_r0 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g2_r1 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g3_r0 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g3_r1 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g4_r0 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g4_r1 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g5_r0 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g5_r1 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g6_r0 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g6_r1 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g7_r0 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g7_r1 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g8_r0 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g8_r1 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g9_r0 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g9_r1 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
XOuterRing iovss sg13g2_GuardRing_P16000W3852HFF
XInnerRing iovdd sg13g2_GuardRing_N15280W3132HTF
XDGATE gate iovdd dpantenna l=0.64um w=0.3um
.ends sg13g2_Clamp_P10N10D

* sg13g2_GuardRing_N7276W2716HFF
.subckt sg13g2_GuardRing_N7276W2716HFF conn

.ends sg13g2_GuardRing_N7276W2716HFF

* sg13g2_DCNDiode
.subckt sg13g2_DCNDiode anode cathode guard
Xdcdiode[0] anode cathode dantenna l=1.26um w=27.78um
Xdcdiode[1] anode cathode dantenna l=1.26um w=27.78um
Xguard guard sg13g2_GuardRing_N7276W2716HFF
.ends sg13g2_DCNDiode

* sg13g2_GuardRing_P7276W2716HFF
.subckt sg13g2_GuardRing_P7276W2716HFF conn

.ends sg13g2_GuardRing_P7276W2716HFF

* sg13g2_DCPDiode
.subckt sg13g2_DCPDiode anode cathode guard
Xdcdiode[0] anode cathode dpantenna l=1.26um w=27.78um
Xdcdiode[1] anode cathode dpantenna l=1.26um w=27.78um
Xguard guard sg13g2_GuardRing_P7276W2716HFF
.ends sg13g2_DCPDiode

* sg13g2_LevelUpInv
.subckt sg13g2_LevelUpInv vdd iovdd vss i o
Xn_i_inv i_n i vss vss sg13_lv_nmos l=0.13um w=2.75um
Xp_i_inv i_n i vdd vdd sg13_lv_pmos l=0.13um w=4.75um
Xn_lvld_n vss i_n lvld_n vss sg13_hv_nmos l=0.45um w=1.9um
Xn_lvld lvld i vss vss sg13_hv_nmos l=0.45um w=1.9um
Xp_lvld_n iovdd lvld lvld_n iovdd sg13_hv_pmos l=0.45um w=0.3um
Xp_lvld lvld lvld_n iovdd iovdd sg13_hv_pmos l=0.45um w=0.3um
Xn_lvld_n_inv vss lvld_n o vss sg13_hv_nmos l=0.45um w=1.9um
Xp_lvld_n_inv iovdd lvld_n o iovdd sg13_hv_pmos l=0.45um w=3.9um
.ends sg13g2_LevelUpInv

* sg13g2_GateLevelUpInv
.subckt sg13g2_GateLevelUpInv vdd vss iovdd core ngate pgate
Xngate_levelup vdd iovdd vss core ngate sg13g2_LevelUpInv
Xpgate_levelup vdd iovdd vss core pgate sg13g2_LevelUpInv
.ends sg13g2_GateLevelUpInv

* sg13g2_IOPadOut20mA
.subckt sg13g2_IOPadOut20mA vss vdd iovss iovdd c2p pad
Xnclamp iovss iovdd pad ngate sg13g2_Clamp_N10N10D
Xpclamp iovss iovdd pad pgate sg13g2_Clamp_P10N10D
Xdcndiode iovss pad iovdd sg13g2_DCNDiode
Xdcpdiode pad iovdd iovss sg13g2_DCPDiode
Xgatelu vdd vss iovdd c2p ngate pgate sg13g2_GateLevelUpInv
.ends sg13g2_IOPadOut20mA
