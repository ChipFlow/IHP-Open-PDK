* sg13g2_IOPadTriOut12mA hierarchy

* sg13g2_GuardRing_N16000W1980HFF
.subckt sg13g2_GuardRing_N16000W1980HFF conn

.ends sg13g2_GuardRing_N16000W1980HFF

* sg13g2_GuardRing_P15280W1260HFF
.subckt sg13g2_GuardRing_P15280W1260HFF conn

.ends sg13g2_GuardRing_P15280W1260HFF

* sg13g2_Clamp_N6N6D
.subckt sg13g2_Clamp_N6N6D iovss iovdd pad gate
Xclamp_g0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g4 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g5 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
XOuterRing iovdd sg13g2_GuardRing_N16000W1980HFF
XInnerRing iovss sg13g2_GuardRing_P15280W1260HFF
XDGATE iovss gate dantenna l=0.64um w=0.3um
.ends sg13g2_Clamp_N6N6D

* sg13g2_GuardRing_P16000W3852HFF
.subckt sg13g2_GuardRing_P16000W3852HFF conn

.ends sg13g2_GuardRing_P16000W3852HFF

* sg13g2_GuardRing_N15280W3132HTF
.subckt sg13g2_GuardRing_N15280W3132HTF conn

.ends sg13g2_GuardRing_N15280W3132HTF

* sg13g2_Clamp_P6N6D
.subckt sg13g2_Clamp_P6N6D iovss iovdd pad gate
Xclamp_g0_r0 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g0_r1 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g1_r0 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g1_r1 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g2_r0 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g2_r1 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g3_r0 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g3_r1 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g4_r0 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g4_r1 iovdd gate pad iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g5_r0 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
Xclamp_g5_r1 pad gate iovdd iovdd sg13_hv_pmos l=0.6um w=6.66um
XOuterRing iovss sg13g2_GuardRing_P16000W3852HFF
XInnerRing iovdd sg13g2_GuardRing_N15280W3132HTF
XDGATE gate iovdd dpantenna l=0.64um w=0.3um
.ends sg13g2_Clamp_P6N6D

* sg13g2_GuardRing_N7276W2716HFF
.subckt sg13g2_GuardRing_N7276W2716HFF conn

.ends sg13g2_GuardRing_N7276W2716HFF

* sg13g2_DCNDiode
.subckt sg13g2_DCNDiode anode cathode guard
Xdcdiode[0] anode cathode dantenna l=1.26um w=27.78um
Xdcdiode[1] anode cathode dantenna l=1.26um w=27.78um
Xguard guard sg13g2_GuardRing_N7276W2716HFF
.ends sg13g2_DCNDiode

* sg13g2_GuardRing_P7276W2716HFF
.subckt sg13g2_GuardRing_P7276W2716HFF conn

.ends sg13g2_GuardRing_P7276W2716HFF

* sg13g2_DCPDiode
.subckt sg13g2_DCPDiode anode cathode guard
Xdcdiode[0] anode cathode dpantenna l=1.26um w=27.78um
Xdcdiode[1] anode cathode dpantenna l=1.26um w=27.78um
Xguard guard sg13g2_GuardRing_P7276W2716HFF
.ends sg13g2_DCPDiode

* tie
.subckt tie vdd vss

.ends tie

* inv_x1
.subckt inv_x1 vdd vss i nq
Xnmos vss i nq vss sg13_lv_nmos l=0.13um w=3.93um
Xpmos vdd i nq vdd sg13_lv_pmos l=0.13um w=4.41um
.ends inv_x1

* nor2_x1
.subckt nor2_x1 vdd vss nq i0 i1
Xi0_nmos vss i0 nq vss sg13_lv_nmos l=0.13um w=3.93um
Xi0_pmos vdd i0 _net0 vdd sg13_lv_pmos l=0.13um w=4.41um
Xi1_nmos nq i1 vss vss sg13_lv_nmos l=0.13um w=3.93um
Xi1_pmos _net0 i1 nq vdd sg13_lv_pmos l=0.13um w=4.41um
.ends nor2_x1

* sg13g2_LevelUp
.subckt sg13g2_LevelUp vdd iovdd vss i o
Xn_i_inv i_n i vss vss sg13_lv_nmos l=0.13um w=2.75um
Xp_i_inv i_n i vdd vdd sg13_lv_pmos l=0.13um w=4.75um
Xn_lvld_n vss i lvld_n vss sg13_hv_nmos l=0.45um w=1.9um
Xn_lvld lvld i_n vss vss sg13_hv_nmos l=0.45um w=1.9um
Xp_lvld_n iovdd lvld lvld_n iovdd sg13_hv_pmos l=0.45um w=0.3um
Xp_lvld lvld lvld_n iovdd iovdd sg13_hv_pmos l=0.45um w=0.3um
Xn_lvld_n_inv vss lvld_n o vss sg13_hv_nmos l=0.45um w=1.9um
Xp_lvld_n_inv iovdd lvld_n o iovdd sg13_hv_pmos l=0.45um w=3.9um
.ends sg13g2_LevelUp

* nand2_x1
.subckt nand2_x1 vdd vss nq i0 i1
Xi0_nmos vss i0 _net0 vss sg13_lv_nmos l=0.13um w=3.93um
Xi0_pmos vdd i0 nq vdd sg13_lv_pmos l=0.13um w=4.41um
Xi1_nmos _net0 i1 nq vss sg13_lv_nmos l=0.13um w=3.93um
Xi1_pmos nq i1 vdd vdd sg13_lv_pmos l=0.13um w=4.41um
.ends nand2_x1

* sg13g2_GateDecode
.subckt sg13g2_GateDecode vdd vss iovdd core en ngate pgate
Xtieinst vdd vss tie
Xen_inv vdd vss en en_n inv_x1
Xngate_nor vdd vss ngate_core core en_n nor2_x1
Xngate_levelup vdd iovdd vss ngate_core ngate sg13g2_LevelUp
Xpgate_nand vdd vss pgate_core core en nand2_x1
Xpgate_levelup vdd iovdd vss pgate_core pgate sg13g2_LevelUp
.ends sg13g2_GateDecode

* sg13g2_IOPadTriOut12mA
.subckt sg13g2_IOPadTriOut12mA vss vdd iovss iovdd c2p c2p_en pad
Xnclamp iovss iovdd pad ngate sg13g2_Clamp_N6N6D
Xpclamp iovss iovdd pad pgate sg13g2_Clamp_P6N6D
Xdcndiode iovss pad iovdd sg13g2_DCNDiode
Xdcpdiode pad iovdd iovss sg13g2_DCPDiode
Xgatedec vdd vss iovdd c2p c2p_en ngate pgate sg13g2_GateDecode
.ends sg13g2_IOPadTriOut12mA
