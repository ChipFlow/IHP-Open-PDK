* sg13g2_IOPadVdd hierarchy

* sg13g2_GuardRing_N16000W4884HFF
.subckt sg13g2_GuardRing_N16000W4884HFF conn

.ends sg13g2_GuardRing_N16000W4884HFF

* sg13g2_GuardRing_P15280W4164HFF
.subckt sg13g2_GuardRing_P15280W4164HFF conn

.ends sg13g2_GuardRing_P15280W4164HFF

* sg13g2_Clamp_N43N43D4R
.subckt sg13g2_Clamp_N43N43D4R iovss iovdd pad gate
Xclamp_g0_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g0_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g0_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g0_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g1_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g1_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g1_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g1_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g2_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g2_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g2_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g2_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g3_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g3_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g3_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g3_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g4_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g4_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g4_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g4_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g5_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g5_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g5_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g5_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g6_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g6_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g6_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g6_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g7_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g7_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g7_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g7_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g8_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g8_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g8_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g8_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g9_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g9_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g9_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g9_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g10_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g10_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g10_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g10_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g11_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g11_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g11_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g11_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g12_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g12_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g12_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g12_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g13_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g13_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g13_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g13_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g14_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g14_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g14_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g14_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g15_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g15_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g15_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g15_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g16_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g16_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g16_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g16_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g17_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g17_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g17_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g17_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g18_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g18_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g18_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g18_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g19_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g19_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g19_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g19_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g20_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g20_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g20_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g20_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g21_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g21_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g21_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g21_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g22_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g22_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g22_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g22_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g23_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g23_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g23_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g23_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g24_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g24_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g24_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g24_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g25_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g25_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g25_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g25_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g26_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g26_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g26_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g26_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g27_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g27_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g27_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g27_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g28_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g28_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g28_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g28_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g29_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g29_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g29_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g29_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g30_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g30_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g30_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g30_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g31_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g31_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g31_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g31_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g32_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g32_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g32_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g32_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g33_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g33_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g33_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g33_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g34_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g34_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g34_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g34_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g35_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g35_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g35_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g35_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g36_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g36_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g36_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g36_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g37_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g37_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g37_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g37_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g38_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g38_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g38_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g38_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g39_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g39_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g39_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g39_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g40_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g40_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g40_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g40_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g41_r0 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g41_r1 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g41_r2 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g41_r3 pad gate iovss iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g42_r0 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g42_r1 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g42_r2 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
Xclamp_g42_r3 iovss gate pad iovss sg13_hv_nmos l=0.6um w=4.4um
XOuterRing iovdd sg13g2_GuardRing_N16000W4884HFF
XInnerRing iovss sg13g2_GuardRing_P15280W4164HFF
XDGATE iovss gate dantenna l=0.64um w=0.3um
.ends sg13g2_Clamp_N43N43D4R

* sg13g2_RCClampResistor
.subckt sg13g2_RCClampResistor pin1 pin2
Rres_fing[0] pin1 conn_0_1 5200.0
Rres_fing[1] conn_0_1 conn_1_2 5200.0
Rres_fing[2] conn_1_2 conn_2_3 5200.0
Rres_fing[3] conn_2_3 conn_3_4 5200.0
Rres_fing[4] conn_3_4 conn_4_5 5200.0
Rres_fing[5] conn_4_5 conn_5_6 5200.0
Rres_fing[6] conn_5_6 conn_6_7 5200.0
Rres_fing[7] conn_6_7 conn_7_8 5200.0
Rres_fing[8] conn_7_8 conn_8_9 5200.0
Rres_fing[9] conn_8_9 conn_9_10 5200.0
Rres_fing[10] conn_9_10 conn_10_11 5200.0
Rres_fing[11] conn_10_11 conn_11_12 5200.0
Rres_fing[12] conn_11_12 conn_12_13 5200.0
Rres_fing[13] conn_12_13 conn_13_14 5200.0
Rres_fing[14] conn_13_14 conn_14_15 5200.0
Rres_fing[15] conn_14_15 conn_15_16 5200.0
Rres_fing[16] conn_15_16 conn_16_17 5200.0
Rres_fing[17] conn_16_17 conn_17_18 5200.0
Rres_fing[18] conn_17_18 conn_18_19 5200.0
Rres_fing[19] conn_18_19 conn_19_20 5200.0
Rres_fing[20] conn_19_20 conn_20_21 5200.0
Rres_fing[21] conn_20_21 conn_21_22 5200.0
Rres_fing[22] conn_21_22 conn_22_23 5200.0
Rres_fing[23] conn_22_23 conn_23_24 5200.0
Rres_fing[24] conn_23_24 conn_24_25 5200.0
Rres_fing[25] conn_24_25 pin2 5200.0
.ends sg13g2_RCClampResistor

* sg13g2_GuardRing_P16000W4466HFT
.subckt sg13g2_GuardRing_P16000W4466HFT conn

.ends sg13g2_GuardRing_P16000W4466HFT

* sg13g2_GuardRing_N9472W2216HTT
.subckt sg13g2_GuardRing_N9472W2216HTT conn

.ends sg13g2_GuardRing_N9472W2216HTT

* sg13g2_RCClampInverter
.subckt sg13g2_RCClampInverter supply ground in out
Xcapmos0_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos1_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos2_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos3_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos4_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos5_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos6_r0 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xnmos0_r0 ground in out ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos1_r0 out in ground ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos2_r0 ground in out ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos3_r0 out in ground ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos4_r0 ground in out ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos5_r0 out in ground ground sg13_hv_nmos l=0.5um w=9.0um
Xcapmos0_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos1_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos2_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos3_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos4_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos5_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xcapmos6_r1 ground in ground ground sg13_hv_nmos l=9.5um w=9.0um
Xnmos0_r1 ground in out ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos1_r1 out in ground ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos2_r1 ground in out ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos3_r1 out in ground ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos4_r1 ground in out ground sg13_hv_nmos l=0.5um w=9.0um
Xnmos5_r1 out in ground ground sg13_hv_nmos l=0.5um w=9.0um
Xnmosguardring ground sg13g2_GuardRing_P16000W4466HFT
Xpmos0_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos1_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos2_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos3_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos4_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos5_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos6_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos7_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos8_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos9_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos10_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos11_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos12_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos13_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos14_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos15_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos16_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos17_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos18_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos19_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos20_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos21_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos22_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos23_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos24_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos25_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos26_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos27_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos28_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos29_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos30_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos31_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos32_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos33_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos34_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos35_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos36_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos37_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos38_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos39_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos40_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos41_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos42_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos43_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos44_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos45_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos46_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos47_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos48_r0 supply in out supply sg13_hv_pmos l=0.5um w=7.0um
Xpmos49_r0 out in supply supply sg13_hv_pmos l=0.5um w=7.0um
Xpmosguardring supply sg13g2_GuardRing_N9472W2216HTT
.ends sg13g2_RCClampInverter

* sg13g2_GuardRing_N7276W2716HFF
.subckt sg13g2_GuardRing_N7276W2716HFF conn

.ends sg13g2_GuardRing_N7276W2716HFF

* sg13g2_DCNDiode
.subckt sg13g2_DCNDiode anode cathode guard
Xdcdiode[0] anode cathode dantenna l=1.26um w=27.78um
Xdcdiode[1] anode cathode dantenna l=1.26um w=27.78um
Xguard guard sg13g2_GuardRing_N7276W2716HFF
.ends sg13g2_DCNDiode

* sg13g2_GuardRing_P7276W2716HFF
.subckt sg13g2_GuardRing_P7276W2716HFF conn

.ends sg13g2_GuardRing_P7276W2716HFF

* sg13g2_DCPDiode
.subckt sg13g2_DCPDiode anode cathode guard
Xdcdiode[0] anode cathode dpantenna l=1.26um w=27.78um
Xdcdiode[1] anode cathode dpantenna l=1.26um w=27.78um
Xguard guard sg13g2_GuardRing_P7276W2716HFF
.ends sg13g2_DCPDiode

* sg13g2_IOPadVdd
.subckt sg13g2_IOPadVdd vss vdd iovss iovdd
Xnclamp iovss iovdd vdd ngate sg13g2_Clamp_N43N43D4R
Xrcres vdd res_cap sg13g2_RCClampResistor
Xrcinv vdd iovss res_cap ngate sg13g2_RCClampInverter
Xdcndiode iovss vdd iovdd sg13g2_DCNDiode
Xdcpdiode vdd iovdd iovss sg13g2_DCPDiode
.ends sg13g2_IOPadVdd
